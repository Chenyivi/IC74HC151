library verilog;
use verilog.vl_types.all;
entity IC74HC151_tb is
end IC74HC151_tb;
