library verilog;
use verilog.vl_types.all;
entity IC74HC151_vlg_vec_tst is
end IC74HC151_vlg_vec_tst;
