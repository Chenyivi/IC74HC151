library verilog;
use verilog.vl_types.all;
entity IC74HC151_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        YF              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end IC74HC151_vlg_check_tst;
